MOS NOR Gate
CL 3 0 .25p

M1 3 1 0 0 NMOD L=3u W=3u
M2 4 1 3 4 PMOD L=3u W=3u
M3 3 2 0 0 NMOD L=3u W=3u
M4 5 2 4 5 PMOD L=3u W=3u

VDD 5 0 DC 5V
VG1 1 0 PULSE(0 5 0 1n 1n 100n 1.5e-7)
VG2 2 0 PULSE(0 0 0 1n 1n 100n 1.5e-7)

.model NMOD NMOS (Level=1 VTO=1 TOX=1e-7)
.model PMOD PMOS (Level=1 VTO=-1 TOX=1e-7)

.control

tran 2e-10 1.5e-7
plot v(1)
plot v(2)
plot v(3)
plot v(4)

.endc

.end
